/*
* File: QUEUE_obj.v
* Author: Nikita Kim & Celine Wang
* Email: kimn1944@gmail.com
* Date: 12/7/19
*/

`include "config.v"

module ROB
    #()
    (input clk,
      input reset,
      input stall,
      input flush,

      input enque,
      input enque_data,

      input deque,

      output deque_data);


endmodule
