


`define LOG_PHYS    $clog2(NUM_PHYS_REGS)

module PhysRegFile #(
    parameter NUM_PHYS_REGS = 64 
)
(
    /* Write Me */
    );
	 
	reg [31:0] PReg [NUM_PHYS_REGS-1:0] /*verilator public*/;

    /* Write Me */
    
endmodule
