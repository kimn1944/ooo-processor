

`define LOG_PHYS    $clog2(NUM_PHYS_REGS)

module RegRead#(
    parameter NUM_PHYS_REGS = 64 
)
(

    /* Write Me */

    );

	PhysRegFile  #(
	.NUM_PHYS_REGS(NUM_PHYS_REGS)
	)
	PhysRegFile(
    /* Write Me */
    );
    
    /* Write Me */
    
endmodule
